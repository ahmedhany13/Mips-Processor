module data_Memory(addr , wdata , rdata , regwrite , regread );

output [31:0] rdata;
input  [31:0] addr;
input  [31:0] wdata;
input  regread;
input  regwrite;

if()



endmodule
